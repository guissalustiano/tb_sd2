-- TODO fix cases of op 1100
-- TODO fix cases of op 0111 (still with SLT values, except for the first)
entity alu_tb is 
end entity;

architecture arch of alu_tb is

    function to_bstring(b : bit) return string is
        variable b_str_v : string(1 to 3);  -- bit image with quotes around
    begin
        b_str_v := bit'image(b);
        return "" & b_str_v(2);  -- "" & character to get string
    end function;

    function to_bstring(bv : bit_vector) return string is
        alias    bv_norm : bit_vector(1 to bv'length) is bv;
        variable b_str_v : string(1 to 1);  -- String of bit
        variable res_v   : string(1 to bv'length);
    begin
        for idx in bv_norm'range loop
            b_str_v := to_bstring(bv_norm(idx));
            res_v(idx) := b_str_v(1);
        end loop;
        return res_v;
    end function;

    component alu is
        generic(
            size: natural := 10
        );
        port(
            A, B: in bit_vector(size-1 downto 0);
            F: out bit_vector(size-1 downto 0);
            S: in bit_vector(3 downto 0);
            Z, Ov, Co: out bit
        );
    end component;

    constant INPUT_SIZE: natural := 10;
    type test_case_type is record
        A: bit_vector(INPUT_SIZE-1 downto 0);
        B: bit_vector(INPUT_SIZE-1 downto 0);
        op: bit_vector(3 downto 0);
        response: bit_vector(INPUT_SIZE-1 downto 0);
    end record;
    type test_case_array is array(1 to 6*INPUT_SIZE) of test_case_type;
    constant TEST_CASES: test_case_array := (
        ("0010101100", "0000111110", "0000", "0000101100"),
        ("0010101100", "0000111110", "0001", "0010111110"),
        ("0010101100", "0000111110", "0010", "0011101010"),
        ("0010101100", "0000111110", "0110", "0001101110"),
        ("0010101100", "0000111110", "0111", "0000111110"),
        ("0010101100", "0000111110", "1100", "1101000001"),
        
        
        ("0110010100", "0101000100", "0000", "0100000100"),
        ("0110010100", "0101000100", "0001", "0111010100"),
        ("0110010100", "0101000100", "0010", "1011011000"),
        ("0110010100", "0101000100", "0110", "0001010000"),
        ("0110010100", "0101000100", "0111", "0101000100"),
        ("0110010100", "0101000100", "1100", "1000101011"),
        
        
        ("0100010111", "0011000001", "0000", "0000000001"),
        ("0100010111", "0011000001", "0001", "0111010111"),
        ("0100010111", "0011000001", "0010", "0111011000"),
        ("0100010111", "0011000001", "0110", "0001010110"),
        ("0100010111", "0011000001", "0111", "0011000001"),
        ("0100010111", "0011000001", "1100", "1000101000"),
        
        
        ("0110101000", "0110001000", "0000", "0110001000"),
        ("0110101000", "0110001000", "0001", "0110101000"),
        ("0110101000", "0110001000", "0010", "1100110000"),
        ("0110101000", "0110001000", "0110", "0000100000"),
        ("0110101000", "0110001000", "0111", "0110001000"),
        ("0110101000", "0110001000", "1100", "1001010111"),
        
        
        ("0111000110", "0000100010", "0000", "0000000010"),
        ("0111000110", "0000100010", "0001", "0111100110"),
        ("0111000110", "0000100010", "0010", "0111101000"),
        ("0111000110", "0000100010", "0110", "0110100100"),
        ("0111000110", "0000100010", "0111", "0000100010"),
        ("0111000110", "0000100010", "1100", "1000011001"),
        
        
        ("0110001010", "0000001100", "0000", "0000001000"),
        ("0110001010", "0000001100", "0001", "0110001110"),
        ("0110001010", "0000001100", "0010", "0110010110"),
        ("0110001010", "0000001100", "0110", "0101111110"),
        ("0110001010", "0000001100", "0111", "0000001100"),
        ("0110001010", "0000001100", "1100", "1001110001"),
        
        
        ("0001001011", "0001000001", "0000", "0001000001"),
        ("0001001011", "0001000001", "0001", "0001001011"),
        ("0001001011", "0001000001", "0010", "0010001100"),
        ("0001001011", "0001000001", "0110", "0000001010"),
        ("0001001011", "0001000001", "0111", "0001000001"),
        ("0001001011", "0001000001", "1100", "1110110100"),
        
        
        ("0110100001", "0000000110", "0000", "0000000000"),
        ("0110100001", "0000000110", "0001", "0110100111"),
        ("0110100001", "0000000110", "0010", "0110100111"),
        ("0110100001", "0000000110", "0110", "0110011011"),
        ("0110100001", "0000000110", "0111", "0000000110"),
        ("0110100001", "0000000110", "1100", "1001011000"),
        
        
        ("0101110100", "0000110100", "0000", "0000110100"),
        ("0101110100", "0000110100", "0001", "0101110100"),
        ("0101110100", "0000110100", "0010", "0110101000"),
        ("0101110100", "0000110100", "0110", "0101000000"),
        ("0101110100", "0000110100", "0111", "0000110100"),
        ("0101110100", "0000110100", "1100", "1010001011"),
        
        
        ("0001010110", "0000001101", "0000", "0000000100"),
        ("0001010110", "0000001101", "0001", "0001011111"),
        ("0001010110", "0000001101", "0010", "0001100011"),
        ("0001010110", "0000001101", "0110", "0001001001"),
        ("0001010110", "0000001101", "0111", "0000001101"),
        ("0001010110", "0000001101", "1100", "1110100000")
    );

    signal A, B, F: bit_vector(INPUT_SIZE-1 downto 0);
    signal opcode: bit_vector(3 downto 0);
    signal zero, overflow, carryOut: bit;

begin

    dut: alu 
        generic map(INPUT_SIZE)
        port map(
            A, B,
            F,
            opcode,
            zero, overflow, carryOut
        );

    tb: process
        variable expected: bit_vector(INPUT_SIZE-1 downto 0);
    begin
        report "BOT";
        for i in TEST_CASES'range loop
            A <= TEST_CASES(i).A;
            B <= TEST_CASES(i).B;
            opcode <= TEST_CASES(i).op;
            expected := TEST_CASES(i).response;
            wait for 1 ps;
            assert F = expected
            report "Test "&integer'image(i)&" failed. "&
                "Expected "&to_bstring(expected)&" "&
                "but got "&to_bstring(F)
            severity warning;
        end loop;
        report "EOT";
        wait;
    end process;

end architecture arch;